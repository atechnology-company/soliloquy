module main

fn c2v_tooling_smoke() {
    println('c2v tooling smoke test passed')
}

fn main() {
    c2v_tooling_smoke()
}
